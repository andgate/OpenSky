// Automatically generated Verilog-2001
module sky(Sw,Led);
  input [1:0] Sw;
  output [1:0] Led;
  Machine_topEntity Machine_topEntity_inst
  (.x (Sw),.result (Led));
endmodule
